// version  N/A
// last edited  PM
// last edited by 
`timescale 1ns / 1ps
module Program_Counter(




);
    always@(*) begin

    end

endmodule